`define NUM_TESTS 155

static bit [127:0] kat_key_vector [0:NUM_TESTS] = {
            128'h0000_0000_0000_0000_0000_0000_0000_0000,
		    128'h0000_0000_0000_0000_0000_0000_0000_0000,
			128'h0000_0000_0000_0000_0000_0000_0000_0000,
			128'h0000_0000_0000_0000_0000_0000_0000_0000,
			128'h0000_0000_0000_0000_0000_0000_0000_0000,
			128'h0000_0000_0000_0000_0000_0000_0000_0000,
			128'h0000_0000_0000_0000_0000_0000_0000_0000,
			128'h10a58869d74be5a374cf867cfb473859,
			128'hcaea65cdbb75e9169ecd22ebe6e54675,
			128'ha2e2fa9baf7d20822ca9f0542f764a41,
			128'hb6364ac4e1de1e285eaf144a2415f7a0,
			128'h64cf9c7abc50b888af65f49d521944b2,
			128'h47d6742eefcc0465dc96355e851b64d9,
			128'h3eb39790678c56bee34bbcdeccf6cdb5,
			128'h64110a924f0743d500ccadae72c13427,
			128'h18d8126516f8a12ab1a36d9f04d68e51,
			128'hf530357968578480b398a3c251cd1093,
			128'hda84367f325d42d601b4326964802e8e,
			128'he37b1c6aa2846f6fdb413f238b089f23,
			128'h6c002b682483e0cabcc731c253be5674,
			128'h143ae8ed6555aba96110ab58893a8ae1,
			128'hb69418a85332240dc82492353956ae0c,
			128'h71b5c08a1993e1362e4d0ce9b22b78d5,
			128'he234cdca2606b81f29408d5f6da21206,
			128'h13237c49074a3da078dc1d828bb78c6f,
			128'h3071a2a48fe6cbd04f1a129098e308f8,
			128'h90f42ec0f68385f2ffc5dfc03a654dce,
	        128'hfebd9a24d8b65c1c787d50a4ed3619a9,
	        128'h80000000000000000000000000000000,
   	        128'hc0000000000000000000000000000000,
	        128'he0000000000000000000000000000000,
	        128'hf0000000000000000000000000000000,
	        128'hf8000000000000000000000000000000,
	        128'hfc000000000000000000000000000000,
	        128'hfe000000000000000000000000000000,
	        128'hff000000000000000000000000000000,
	        128'hff800000000000000000000000000000,
	        128'hffc00000000000000000000000000000,
	        128'hffe00000000000000000000000000000,
	        128'hfff00000000000000000000000000000,
	        128'hfff80000000000000000000000000000,
	        128'hfffc0000000000000000000000000000,
	        128'hfffe0000000000000000000000000000,
	        128'hffff0000000000000000000000000000,
	        128'hffff8000000000000000000000000000,
	        128'hffffc000000000000000000000000000,
	        128'hffffe000000000000000000000000000,
	        128'hfffff000000000000000000000000000,
	        128'hfffff800000000000000000000000000,
	        128'hfffffc00000000000000000000000000,
	        128'hfffffe00000000000000000000000000,
	        128'hffffff00000000000000000000000000,
	        128'hffffff80000000000000000000000000,
	        128'hffffffc0000000000000000000000000,
	        128'hffffffe0000000000000000000000000,
	        128'hfffffff0000000000000000000000000,
	        128'hfffffff8000000000000000000000000,
	        128'hfffffffc000000000000000000000000,
	        128'hfffffffe000000000000000000000000,
	        128'hffffffff000000000000000000000000,
	        128'hffffffff800000000000000000000000,
	        128'hffffffffc00000000000000000000000,
	        128'hffffffffe00000000000000000000000,
	        128'hfffffffff00000000000000000000000,
	        128'hfffffffff80000000000000000000000,
	        128'hfffffffffc0000000000000000000000,
	        128'hfffffffffe0000000000000000000000,
	        128'hffffffffff0000000000000000000000,
	        128'hffffffffff8000000000000000000000,
	        128'hffffffffffc000000000000000000000,
	        128'hffffffffffe000000000000000000000,
	        128'hfffffffffff000000000000000000000,
	        128'hfffffffffff800000000000000000000,
	        128'hfffffffffffc00000000000000000000,
	        128'hfffffffffffe00000000000000000000,
	        128'hffffffffffff00000000000000000000,
	        128'hffffffffffff80000000000000000000,
	        128'hffffffffffffc0000000000000000000,
	        128'hffffffffffffe0000000000000000000,
	        128'hfffffffffffff0000000000000000000,
	        128'hfffffffffffff8000000000000000000,
	        128'hfffffffffffffc000000000000000000,
	        128'hfffffffffffffe000000000000000000,
	        128'hffffffffffffff000000000000000000,
	        128'hffffffffffffff800000000000000000,
	        128'hffffffffffffffc00000000000000000,
	        128'hffffffffffffffe00000000000000000,
	        128'hfffffffffffffff00000000000000000,
	        128'hfffffffffffffff80000000000000000,
	        128'hfffffffffffffffc0000000000000000,
	        128'hfffffffffffffffe0000000000000000,
	        128'hffffffffffffffff0000000000000000,
	        128'hffffffffffffffff8000000000000000,
	        128'hffffffffffffffffc000000000000000,
	        128'hffffffffffffffffe000000000000000,
	        128'hfffffffffffffffff000000000000000,
	        128'hfffffffffffffffff800000000000000,
	        128'hfffffffffffffffffc00000000000000,
	        128'hfffffffffffffffffe00000000000000,
	        128'hffffffffffffffffff00000000000000,
	        128'hffffffffffffffffff80000000000000,
	        128'hffffffffffffffffffc0000000000000,
	        128'hffffffffffffffffffe0000000000000,
	        128'hfffffffffffffffffff0000000000000,
	        128'hfffffffffffffffffff8000000000000,
	        128'hfffffffffffffffffffc000000000000,
	        128'hfffffffffffffffffffe000000000000,
	        128'hffffffffffffffffffff000000000000,
	        128'hffffffffffffffffffff800000000000,
	        128'hffffffffffffffffffffc00000000000,
	        128'hffffffffffffffffffffe00000000000,
	        128'hfffffffffffffffffffff00000000000,
	        128'hfffffffffffffffffffff80000000000,
	        128'hfffffffffffffffffffffc0000000000,
	        128'hfffffffffffffffffffffe0000000000,
	        128'hffffffffffffffffffffff0000000000,
	        128'hffffffffffffffffffffff8000000000,
	        128'hffffffffffffffffffffffc000000000,
	        128'hffffffffffffffffffffffe000000000,
	        128'hfffffffffffffffffffffff000000000,
	        128'hfffffffffffffffffffffff800000000,
	        128'hfffffffffffffffffffffffc00000000,
	        128'hfffffffffffffffffffffffe00000000,
	        128'hffffffffffffffffffffffff00000000,
	        128'hffffffffffffffffffffffff80000000,
	        128'hffffffffffffffffffffffffc0000000,
	        128'hffffffffffffffffffffffffe0000000,
	        128'hfffffffffffffffffffffffff0000000,
	        128'hfffffffffffffffffffffffff8000000,
	        128'hfffffffffffffffffffffffffc000000,
	        128'hfffffffffffffffffffffffffe000000,
	        128'hffffffffffffffffffffffffff000000,
	        128'hffffffffffffffffffffffffff800000,
	        128'hffffffffffffffffffffffffffc00000,
	        128'hffffffffffffffffffffffffffe00000,
	        128'hfffffffffffffffffffffffffff00000,
	        128'hfffffffffffffffffffffffffff80000,
	        128'hfffffffffffffffffffffffffffc0000,
	        128'hfffffffffffffffffffffffffffe0000,
	        128'hffffffffffffffffffffffffffff0000,
	        128'hffffffffffffffffffffffffffff8000,
	        128'hffffffffffffffffffffffffffffc000,
	        128'hffffffffffffffffffffffffffffe000,
	        128'hfffffffffffffffffffffffffffff000,
	        128'hfffffffffffffffffffffffffffff800,
	        128'hfffffffffffffffffffffffffffffc00,
	        128'hfffffffffffffffffffffffffffffe00,
	        128'hffffffffffffffffffffffffffffff00,
	        128'hffffffffffffffffffffffffffffff80,
	        128'hffffffffffffffffffffffffffffffc0,
	        128'hffffffffffffffffffffffffffffffe0,
	        128'hfffffffffffffffffffffffffffffff0,
	        128'hfffffffffffffffffffffffffffffff8,
	        128'hfffffffffffffffffffffffffffffffc,
	        128'hfffffffffffffffffffffffffffffffe,
	        128'hffffffffffffffffffffffffffffffff};
					     

static bit [127:0] kat_plain_vector [0:NUM_TESTS] = {
           128'hf344_81ec_3cc6_27ba_cd5d_c3fb_08f2_73e6,
		   128'h9798_c464_0bad_75c7_c322_7db9_1017_4e72,
		   128'h96ab_5c2f_f612_d9df_aae8_c31f_30c4_2168,
		   128'h6a11_8a87_4519_e64e_9963_798a_503f_1d35,
		   128'hcb9f_ceec_8128_6ca3_e989_bd97_9b0c_b284,
		   128'hb26a_eb18_74e4_7ca8_358f_f223_78f0_9144,
		   128'h58c8_e00b_2631_686d_54ea_b84b_91f0_aca1,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000,
		   128'h00000000000000000000000000000000};
		   

static bit [127:0] kat_cipher_vector [0:NUM_TESTS] = {
            128'h0336_763e_966d_9259_5a56_7cc9_ce53_7f5e,
		    128'ha9a1_631b_f499_6954_ebc0_9395_7b23_4589,
		    128'hff4f_8391_a6a4_0ca5_b25d_23be_dd44_a597,
		    128'hdc43_be40_be0e_5371_2f7e_2bf5_ca70_7209,
		    128'h92be_edab_1895_a94f_aa69_b632_e5cc_47ce,
		    128'h4592_64f4_798f_6a78_bacb_89c1_5ed3_d601,
		    128'h08a4_e2ef_ec8a_8e33_12ca_7460_b904_0bbf,
		    128'h6d251e6944b051e04eaa6fb4dbf78465,
		    128'h6e29201190152df4ee058139def610bb,
		    128'hc3b44b95d9d2f25670eee9a0de099fa3,
		    128'h5d9b05578fc944b3cf1ccf0e746cd581,
		    128'hf7efc89d5dba578104016ce5ad659c05,
		    128'h0306194f666d183624aa230a8b264ae7,
		    128'h858075d536d79ccee571f7d7204b1f67,
			128'h35870c6a57e9e92314bcb8087cde72ce,
			128'h6c68e9be5ec41e22c825b7c7affb4363,
			128'hf5df39990fc688f1b07224cc03e86cea,
			128'hbba071bcb470f8f6586e5d3add18bc66,
			128'h43c9f7e62f5d288bb27aa40ef8fe1ea8,
			128'h3580d19cff44f1014a7c966a69059de5,
			128'h806da864dd29d48deafbe764f8202aef,
			128'ha303d940ded8f0baff6f75414cac5243,
			128'hc2dabd117f8a3ecabfbb11d12194d9d0,
			128'hfff60a4740086b3b9c56195b98d91a7b,
			128'h8146a08e2357f0caa30ca8c94d1a0544,
			128'h4b98e06d356deb07ebb824e5713f7be3,
			128'h7a20a53d460fc9ce0423a7a0764c6cf2,
			128'hf4a70d8af877f9b02b4c40df57d45b17,
			128'h0edd33d3c621e546455bd8ba1418bec8,
			128'h4bc3f883450c113c64ca42e1112a9e87,
			128'h72a1da770f5d7ac4c9ef94d822affd97,
			128'h970014d634e2b7650777e8e84d03ccd8,
			128'hf17e79aed0db7e279e955b5f493875a7,
			128'h9ed5a75136a940d0963da379db4af26a,
			128'hc4295f83465c7755e8fa364bac6a7ea5,
			128'hb1d758256b28fd850ad4944208cf1155,
			128'h42ffb34c743de4d88ca38011c990890b,
			128'h9958f0ecea8b2172c0c1995f9182c0f3,
			128'h956d7798fac20f82a8823f984d06f7f5,
			128'ha01bf44f2d16be928ca44aaf7b9b106b,
			128'hb5f1a33e50d40d103764c76bd4c6b6f8,
			128'h2637050c9fc0d4817e2d69de878aee8d,
			128'h113ecbe4a453269a0dd26069467fb5b5,
			128'h97d0754fe68f11b9e375d070a608c884,
			128'hc6a0b3e998d05068a5399778405200b4,
			128'hdf556a33438db87bc41b1752c55e5e49,
			128'h90fb128d3a1af6e548521bb962bf1f05,
			128'h26298e9c1db517c215fadfb7d2a8d691,
			128'ha6cb761d61f8292d0df393a279ad0380,
			128'h12acd89b13cd5f8726e34d44fd486108,
			128'h95b1703fc57ba09fe0c3580febdd7ed4,
			128'hde11722d893e9f9121c381becc1da59a,
			128'h6d114ccb27bf391012e8974c546d9bf2,
			128'h5ce37e17eb4646ecfac29b9cc38d9340,
			128'h18c1b6e2157122056d0243d8a165cddb,
			128'h99693e6a59d1366c74d823562d7e1431,
			128'h6c7c64dc84a8bba758ed17eb025a57e3,
			128'he17bc79f30eaab2fac2cbbe3458d687a,
			128'h1114bc2028009b923f0b01915ce5e7c4,
			128'h9c28524a16a1e1c1452971caa8d13476,
			128'hed62e16363638360fdd6ad62112794f0,
			128'h5a8688f0b2a2c16224c161658ffd4044,
			128'h23f710842b9bb9c32f26648c786807ca,
			128'h44a98bf11e163f632c47ec6a49683a89,
			128'h0f18aff94274696d9b61848bd50ac5e5,
			128'h82408571c3e2424540207f833b6dda69,
			128'h303ff996947f0c7d1f43c8f3027b9b75,
			128'h7df4daf4ad29a3615a9b6ece5c99518a,
			128'hc72954a48d0774db0b4971c526260415,
			128'h1df9b76112dc6531e07d2cfda04411f0,
			128'h8e4d8e699119e1fc87545a647fb1d34f,
			128'he6c4807ae11f36f091c57d9fb68548d1,
			128'h8ebf73aad49c82007f77a5c1ccec6ab4,
			128'h4fb288cc2040049001d2c7585ad123fc,
			128'h04497110efb9dceb13e2b13fb4465564,
			128'h75550e6cb5a88e49634c9ab69eda0430,
			128'hb6768473ce9843ea66a81405dd50b345,
			128'hcb2f430383f9084e03a653571e065de6,
			128'hff4e66c07bae3e79fb7d210847a3b0ba,
			128'h7b90785125505fad59b13c186dd66ce3,
			128'h8b527a6aebdaec9eaef8eda2cb7783e5,
			128'h43fdaf53ebbc9880c228617d6a9b548b,
			128'h53786104b9744b98f052c46f1c850d0b,
			128'hb5ab3013dd1e61df06cbaf34ca2aee78,
			128'h7470469be9723030fdcc73a8cd4fbb10,
			128'ha35a63f5343ebe9ef8167bcb48ad122e,
			128'hfd8687f0757a210e9fdf181204c30863,
			128'h7a181e84bd5457d26a88fbae96018fb0,
			128'h653317b9362b6f9b9e1a580e68d494b5,
			128'h995c9dc0b689f03c45867b5faa5c18d1,
			128'h77a4d96d56dda398b9aabecfc75729fd,
			128'h84be19e053635f09f2665e7bae85b42d,
			128'h32cd652842926aea4aa6137bb2be2b5e,
			128'h493d4a4f38ebb337d10aa84e9171a554,
			128'hd9bff7ff454b0ec5a4a2a69566e2cb84,
			128'h3535d565ace3f31eb249ba2cc6765d7a,
			128'hf60e91fc3269eecf3231c6e9945697c6,
			128'hab69cfadf51f8e604d9cc37182f6635a,
			128'h7866373f24a0b6ed56e0d96fcdafb877,
			128'h1ea448c2aac954f5d812e9d78494446a,
			128'hacc5599dd8ac02239a0fef4a36dd1668,
			128'hd8764468bb103828cf7e1473ce895073,
			128'h1b0d02893683b9f180458e4aa6b73982,
			128'h96d9b017d302df410a937dcdb8bb6e43,
			128'hef1623cc44313cff440b1594a7e21cc6,
			128'h284ca2fa35807b8b0ae4d19e11d7dbd7,
			128'hf2e976875755f9401d54f36e2a23a594,
			128'hec198a18e10e532403b7e20887c8dd80,
			128'h545d50ebd919e4a6949d96ad47e46a80,
			128'hdbdfb527060e0a71009c7bb0c68f1d44,
			128'h9cfa1322ea33da2173a024f2ff0d896d,
			128'h8785b1a75b0f3bd958dcd0e29318c521,
			128'h38f67b9e98e4a97b6df030a9fcdd0104,
			128'h192afffb2c880e82b05926d0fc6c448b,
			128'h6a7980ce7b105cf530952d74daaf798c,
			128'hea3695e1351b9d6858bd958cf513ef6c,
			128'h6da0490ba0ba0343b935681d2cce5ba1,
			128'hf0ea23af08534011c60009ab29ada2f1,
			128'hff13806cf19cc38721554d7c0fcdcd4b,
			128'h6838af1f4f69bae9d85dd188dcdf0688,
			128'h36cf44c92d550bfb1ed28ef583ddf5d7,
			128'hd06e3195b5376f109d5c4ec6c5d62ced,
			128'hc440de014d3d610707279b13242a5c36,
			128'hf0c5c6ffa5e0bd3a94c88f6b6f7c16b9,
			128'h3e40c3901cd7effc22bffc35dee0b4d9,
			128'hb63305c72bedfab97382c406d0c49bc6,
			128'h36bbaab22a6bd4925a99a2b408d2dbae,
			128'h307c5b8fcd0533ab98bc51e27a6ce461,
			128'h829c04ff4c07513c0b3ef05c03e337b5,
			128'hf17af0e895dda5eb98efc68066e84c54,
			128'h277167f3812afff1ffacb4a934379fc3,
			128'h2cb1dc3a9c72972e425ae2ef3eb597cd,
			128'h36aeaa3a213e968d4b5b679d3a2c97fe,
			128'h9241daca4fdd034a82372db50e1a0f3f,
			128'hc14574d9cd00cf2b5a7f77e53cd57885,
			128'h793de39236570aba83ab9b737cb521c9,
			128'h16591c0f27d60e29b85a96c33861a7ef,
			128'h44fb5c4d4f5cb79be5c174a3b1c97348,
			128'h674d2b61633d162be59dde04222f4740,
			128'hb4750ff263a65e1f9e924ccfd98f3e37,
			128'h62d0662d6eaeddedebae7f7ea3a4f6b6,
			128'h70c46bb30692be657f7eaa93ebad9897,
			128'h323994cfb9da285a5d9642e1759b224a,
			128'h1dbf57877b7b17385c85d0b54851e371,
			128'hdfa5c097cdc1532ac071d57b1d28d1bd,
			128'h3a0c53fa37311fc10bd2a9981f513174,
			128'hba4f970c0a25c41814bdae2e506be3b4,
			128'h2dce3acb727cd13ccd76d425ea56e4f6,
			128'h5160474d504b9b3eefb68d35f245f4b3,
			128'h41a8a947766635dec37553d9a6c0cbb7,
			128'h25d6cfe6881f2bf497dd14cd4ddf445b,
			128'h41c78c135ed9e98c096640647265da1e,
			128'h5a4d404d8917e353e92a21072c3b2305,
			128'h02bc96846b3fdc71643f384cd3cc3eaf,
			128'h9ba4a9143f4e5d4048521c4f8877d88e,
			128'ha1f6258c877d5fcd8964484538bfc92c};

